LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;


ENTITY CCR IS
	PORT (
	CLK: IN STD_LOGIC;
	CCR_EN: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	CCR_VALUE: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
	CCR_OUT: OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
	RST: IN STD_LOGIC);
END ENTITY;


ARCHITECTURE CCR_A OF CCR is
COMPONENT onebit_reg
PORT( 
Clk,Rst,En : IN std_logic;
d : IN std_logic_vector(2 DOWNTO 0);
q : OUT std_logic_vector(2 DOWNTO 0));
END COMPONENT;
-----------------------------------------------------
SIGNAL EN, Z, N, C: STD_LOGIC;
SIGNAL FLAG_VALUE, FLAG_READ: STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
BEGIN
EN <= CCR_EN(0) OR CCR_EN(1) OR CCR_EN(2);

Z <=  FLAG_READ(0) WHEN CCR_VALUE(0) = 'Z' OR CCR_EN(0) = '0'
ELSE CCR_VALUE(0) WHEN CCR_EN(0) = '1';

N <=  FLAG_READ(1) WHEN CCR_VALUE(1) = 'Z' OR CCR_EN(1) = '0'
ELSE CCR_VALUE(1) WHEN CCR_EN(1) = '1';

C <=  FLAG_READ(2) WHEN CCR_VALUE(2) = 'Z' OR CCR_EN(2) = '0'
ELSE CCR_VALUE(2) WHEN CCR_EN(2) = '1';

FLAG_VALUE(0)<= Z;
FLAG_VALUE(1)<= N;
FLAG_VALUE(2)<= C;
Flag: onebit_reg PORT MAP(CLK, RST, EN, FLAG_VALUE, FLAG_READ);
CCR_OUT <= FLAG_READ;
END CCR_A;
